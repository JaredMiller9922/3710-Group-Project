// This is the datapath module
module datapath #(paramter REGBITS = 3)
(

	// Create localparams
	
	// Create wires
	
	
	// datapath registers and muxes 
	
	// Instantiate the register file and the alu
);

endmodule 