module GroupProject3710 ();





endmodule